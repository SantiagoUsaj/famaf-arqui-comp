`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.09.2025 11:25:10
// Design Name: 
// Module Name: imem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module imem
    #(parameter N = 32) 
    (
        input logic [6:0] addr, // Agregamos un bit mas para direccionar 128 instrucciones
        output logic [N-1:0] q
    );

    logic [N-1:0] ROM [0:127] = '{default: 32'h0}; // Se agrega espacio para 128 instrucciones

	initial begin
        // Codigo original   
        /*
		ROM [0:46] ='{  32'hf8000001,
                        32'hf8008002,
                        32'hf8000203,
                        32'h8b050083,
                        32'hf8018003,
                        32'hcb050083,
                        32'hf8020003,
                        32'hcb0a03e4,
                        32'hf8028004,
                        32'h8b040064,
                        32'hf8030004,
                        32'hcb030025,
                        32'hf8038005,
                        32'h8a1f0145,
                        32'hf8040005,
                        32'h8a030145,
                        32'hf8048005,
                        32'h8a140294,
                        32'hf8050014,
                        32'haa1f0166,
                        32'hf8058006,
                        32'haa030166,
                        32'hf8060006,
                        32'hf840000c,
                        32'h8b1f0187,
                        32'hf8068007,
                        32'hf807000c,
                        32'h8b0e01bf,
                        32'hf807801f,
                        32'hb4000040,
                        32'hf8080015,
                        32'hf8088015,
                        32'h8b0103e2,
                        32'hcb010042,
                        32'h8b0103f8,
                        32'hf8090018,
                        32'h8b080000,
                        32'hb4ffff82,
                        32'hf809001e,
                        32'h8b1e03de,
                        32'hcb1503f5,
                        32'h8b1403de,
                        32'hf85f83d9,
                        32'h8b1e03de,
                        32'h8b1003de,
                        32'hf81f83d9,
                        32'hb400001f};
        */

        // Codigo modificado para los hazards
              /*
        ROM [0:87] ='{  32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'h8b050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018003,
                        32'hcb050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8020003,
                        32'hcb0a03e4,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8028004,
                        32'h8b040064,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8030004,
                        32'hcb030025,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8038005,
                        32'h8a1f0145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8040005,
                        32'h8a030145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8048005,
                        32'h8a140294,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8050014,
                        32'haa1f0166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8058006,
                        32'haa030166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8060006,
                        32'hf840000c,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f0187,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8068007,
                        32'hf807000c,
                        32'h8b0e01bf,
                        32'hf807801f,
                        32'hb40000a0,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8080015,
                        32'hf8088015,
                        32'h8b0103e2,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb010042,
                        32'h8b0103f8,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8090018,
                        32'h8b080000,
                        32'hb4ffff42,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf809001e,
                        32'h8b1e03de,
                        32'hcb1503f5,
                        32'h8b1f03ff,
                        32'h8b1403de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf85f83d9,
                        32'h8b1e03de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1003de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf81f83d9,
                        32'hb400001f};
        */

        // Codigo con LSL y LSR
        /*
        ROM [0:9] ='{   32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'hd3620884,
                        32'hd34104c6,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018004,
                        32'hf8020006,
                        32'hb400001f};
        */

        // Codigo Juego con LEDS y Switches        
        
        ROM [0:126] ='{
32'h8b0103e6,
32'h8b1f03e0,
32'h8b1f03e1,
32'h8b1f03e2,
32'h8b1f03e3,
32'h8b1f03e4,
32'h8b1f03e5,
32'h8b1f03e7,
32'h8b1f03e8,
32'h8b060000,
32'h8b1f03ff,
32'h8b1f03ff,
32'hd37f3c00,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'hd37f3c21,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b060021,
32'h8b0603e2,
32'h8b1f03e3,
32'h8b0603e4,
32'h8b1f03ff,
32'h8b1f03ff,
32'hd37f0884,
32'h8b0603e7,
32'h8b1f03ff,
32'h8b1f03ff,
32'hd37f3ce7,
32'h8b0603e8,
32'hf8000002,
32'hf8400025,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8a0600a5,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb4000125,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b0603e3,
32'hb40000ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03e3,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb40002e3,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hd35f0442,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8a08004a,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb400012a,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b0703e2,
32'hb400037f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb40002ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hd37f0442,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8a07004a,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb400012a,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b0803e2,
32'hb400011f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb400009f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b0403e9,
32'h8b1f03ff,
32'h8b1f03ff,
32'hcb060129,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb4fff7a9,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb4ffff3f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff};

         
	end

	always_comb begin
		q = ROM[addr];
	end

endmodule


