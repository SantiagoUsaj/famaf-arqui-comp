`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.09.2025 11:25:10
// Design Name: 
// Module Name: imem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module imem
    #(parameter N = 32) 
    (
        input logic [6:0] addr, // Agregamos un bit mas para direccionar 128 instrucciones
        output logic [N-1:0] q
    );

    logic [N-1:0] ROM [0:127] = '{default: 32'h0}; // Se agrega espacio para 128 instrucciones

	initial begin      

        // Codigo original modificado con NOPS
        /*
        ROM [0:87] ='{  32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'h8b050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018003,
                        32'hcb050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8020003,
                        32'hcb0a03e4,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8028004,
                        32'h8b040064,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8030004,
                        32'hcb030025,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8038005,
                        32'h8a1f0145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8040005,
                        32'h8a030145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8048005,
                        32'h8a140294,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8050014,
                        32'haa1f0166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8058006,
                        32'haa030166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8060006,
                        32'hf840000c,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f0187,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8068007,
                        32'hf807000c,
                        32'h8b0e01bf,
                        32'hf807801f,
                        32'hb40000a0,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8080015,
                        32'hf8088015,
                        32'h8b0103e2,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb010042,
                        32'h8b0103f8,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8090018,
                        32'h8b080000,
                        32'hb4ffff42,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf809001e,
                        32'h8b1e03de,
                        32'hcb1503f5,
                        32'h8b1f03ff,
                        32'h8b1403de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf85f83d9,
                        32'h8b1e03de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1003de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf81f83d9,
                        32'hb400001f};
        */
        
        // Codigo base para probar el funcionamiento de LSL y LSR
        /*
        ROM [0:9] ='{   32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'hd3620884,
                        32'hd34104c6,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018004,
                        32'hf8020006,
                        32'hb400001f
                    };
        */

        // Codigo original modificado con NOPS , LSL y LSR
        ROM [0:87] ='{  32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'h8b050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018003,
                        32'hcb050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8020003,
                        32'hcb0a03e4,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8028004,
                        32'h8b040064,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8030004,
                        32'hcb030025,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8038005,
                        32'h8a1f0145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8040005,
                        32'h8a030145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8048005,
                        32'h8a140294,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8050014,
                        32'hd35f0966,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8058006,
                        32'haa030166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8060006,
                        32'hf840000c,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f1187,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8068007,
                        32'hf807000c,
                        32'h8b0e01bf,
                        32'hf807801f,
                        32'hb40000a0,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8080015,
                        32'hf8088015,
                        32'h8b0103e2,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb010042,
                        32'h8b0103f8,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8090018,
                        32'h8b080000,
                        32'hb4ffff42,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf809001e,
                        32'h8b1e03de,
                        32'hcb1503f5,
                        32'h8b1f03ff,
                        32'h8b1403de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf85f83d9,
                        32'h8b1e03de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1003de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf81f83d9,
                        32'hb400001f};
            
         // Leds con sw0 y sw1
         /*
         ROM [0:103] ='{
                            32'h8b0103ea,
                            32'h8b0203eb,
                            32'h8b0103e4,
                            32'h8b1f03e0,
                            32'h8b1f03e1,
                            32'h8b1f03e2,
                            32'h8b1f03e3,
                            32'h8b1f03e5,
                            32'h8b040000,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f3c00,
                            32'h8b040021,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f3c21,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b080021,
                            32'h8b0403e3,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f4063,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hcb040063,
                            32'h8b0403e5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'hf8400022,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8a0a0054,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4000114,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hf8000003,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4fffe7f,
                            32'h8a0b0055,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4000175,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hf8000005,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4fffd1f,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hf800001f,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4fffc3f,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff};
        */
	end
	always_comb begin
		q = ROM[addr];
	end

endmodule


