`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.09.2025 09:53:16
// Design Name: 
// Module Name: mux2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2 
    #(parameter N = 64)
    (
        input logic [N-1:0] d0, d1,
        input logic s,
        output logic [N-1:0] y
    );
				
	assign y = s ? d1 : d0;
	
endmodule

