`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.09.2025 11:25:10
// Design Name: 
// Module Name: imem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module imem
    #(parameter N = 32) 
    (
        input logic [5:0] addr, // Agregamos 1 bit mas para direccionar 128 instrucciones - Luego se cambio a 8 bits para direccionar 256 instrucciones por los leds y switches
        output logic [N-1:0] q
    );

    logic [N-1:0] ROM [0:63] = '{default: 32'h0}; // Se agrega espacio para 128 instrucciones - Luego se cambio a 256 instrucciones para los leds y switches

	initial begin      

        // original_code_nops.s
        /*
        ROM [0:87] ='{  32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'h8b050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018003,
                        32'hcb050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8020003,
                        32'hcb0a03e4,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8028004,
                        32'h8b040064,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8030004,
                        32'hcb030025,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8038005,
                        32'h8a1f0145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8040005,
                        32'h8a030145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8048005,
                        32'h8a140294,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8050014,
                        32'haa1f0166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8058006,
                        32'haa030166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8060006,
                        32'hf840000c,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f0187,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8068007,
                        32'hf807000c,
                        32'h8b0e01bf,
                        32'hf807801f,
                        32'hb40000a0,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8080015,
                        32'hf8088015,
                        32'h8b0103e2,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb010042,
                        32'h8b0103f8,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8090018,
                        32'h8b080000,
                        32'hb4ffff42,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf809001e,
                        32'h8b1e03de,
                        32'hcb1503f5,
                        32'h8b1f03ff,
                        32'h8b1403de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf85f83d9,
                        32'h8b1e03de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1003de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf81f83d9,
                        32'hb400001f};
        */
        
        // basic_shift.s
        /*
        ROM [0:9] ='{   32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'hd3620884,
                        32'hd34104c6,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018004,
                        32'hf8020006,
                        32'hb400001f
                    };
        */

        // original_code_nops_ls.s
        /*
        ROM [0:87] ='{  32'hf8000001,
                        32'hf8008002,
                        32'hf8010003,
                        32'h8b050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8018003,
                        32'hcb050083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8020003,
                        32'hcb0a03e4,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8028004,
                        32'h8b040064,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8030004,
                        32'hcb030025,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8038005,
                        32'h8a1f0145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8040005,
                        32'h8a030145,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8048005,
                        32'h8a140294,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8050014,
                        32'hd35f0966,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8058006,
                        32'haa030166,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8060006,
                        32'hf840000c,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f1187,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8068007,
                        32'hf807000c,
                        32'h8b0e01bf,
                        32'hf807801f,
                        32'hb40000a0,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8080015,
                        32'hf8088015,
                        32'h8b0103e2,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb010042,
                        32'h8b0103f8,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8090018,
                        32'h8b080000,
                        32'hb4ffff42,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf809001e,
                        32'h8b1e03de,
                        32'hcb1503f5,
                        32'h8b1f03ff,
                        32'h8b1403de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf85f83d9,
                        32'h8b1e03de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1003de,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf81f83d9,
                        32'hb400001f};
            */
            
         // off_on_even.s
         /*
         ROM [0:103] ='{
                            32'h8b0103ea,
                            32'h8b0203eb,
                            32'h8b0103e4,
                            32'h8b1f03e0,
                            32'h8b1f03e1,
                            32'h8b1f03e2,
                            32'h8b1f03e3,
                            32'h8b1f03e5,
                            32'h8b040000,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f3c00,
                            32'h8b040021,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f3c21,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b080021,
                            32'h8b0403e3,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f4063,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hcb040063,
                            32'h8b0403e5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hd37f08a5,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b0400a5,
                            32'hf8400022,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8a0a0054,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4000114,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hf8000003,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4fffe7f,
                            32'h8a0b0055,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4000175,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hf8000005,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4fffd1f,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hf800001f,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'hb4fffc3f,
                            32'h8b1f03ff,
                            32'h8b1f03ff,
                            32'h8b1f03ff};
        */
        // expansion.s
        /*
       ROM [0:114] ='{
                        32'h8b0103e4,
                        32'h8b1f03e0,
                        32'h8b1f03e1,
                        32'h8b1f03e2,
                        32'h8b1f03e3,
                        32'h8b1f03e5,
                        32'h8b1f03e6,
                        32'h8b1f03ea,
                        32'h8b1f03eb,
                        32'h8b040000,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f3c00,
                        32'h8b040021,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f3c21,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b080021,
                        32'h8b0403e5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'hd37f0483,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b040063,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f1c63,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f006b,
                        32'hf8000003,
                        32'h8b0503ea,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb04014a,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb400010a,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4ffff3f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8400022,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8a040042,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000162,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0b03e3,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4fffc9f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f0467,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd35f0468,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'haa070063,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'haa080063,
                        32'hd37f4086,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb0400c6,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb060067,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000107,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4fff93f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8000003,
                        32'h8b0503ea,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb04014a,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb400010a,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4ffff3f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0b03e3,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4fff67f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff};
        */
	/*
        // leds_and_switches.s
        ROM [0:187] ='{
                        32'h8b0103e4,
                        32'h8b0203ec,
                        32'h8b0403ed,
                        32'h8b1f03e0,
                        32'h8b1f03e1,
                        32'h8b1f03e2,
                        32'h8b1f03e3,
                        32'h8b1f03e5,
                        32'h8b1f03e6,
                        32'h8b1f03e7,
                        32'h8b1f03e9,
                        32'h8b1f03ea,
                        32'h8b1f03eb,
                        32'hd37f3c80,
                        32'hd37f3c81,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b080021,
                        32'hd37f4083,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb040063,
                        32'hd37f0885,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f08a5,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0400a5,
                        32'hd37f088a,
                        32'hd37f048b,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b04016b,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f1d6b,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8400022,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8a040046,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000126,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8000003,
                        32'hb4fffebf,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8a0c0046,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000126,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8000005,
                        32'hb4fffd3f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8a0d0046,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000a26,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0b03e8,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8000008,
                        32'h8b0a03e9,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb040129,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000109,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4ffff3f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8400022,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8a040046,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000106,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4fff85f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f0507,
                        32'hd35f0509,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'haa070108,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'haa090108,
                        32'hd37f4086,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb0400c6,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb060107,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000107,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4fff9df,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8000008,
                        32'h8b0a03e9,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb040129,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4000109,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb4ffff3f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b0b03e8,
                        32'hb4fff75f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf800001f,
                        32'hb4fff21f,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'h8b1f03ff
                    };
                    */

        // solo prender leds
        /*
        ROM [0:21] ='{
                        32'h8b0103e4,
                        32'h8b1f03e0,
                        32'h8b1f03e1,
                        32'h8b1f03e2,
                        32'h8b1f03e3,
                        32'h8b040000,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f3c00,
                        32'h8b0403e3,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hd37f4063,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hcb040063,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hf8000003,
                        32'h8b1f03ff,
                        32'h8b1f03ff,
                        32'hb400001f};
                        */
    ROM [0:30] ='{
                    32'h8b0103e4,
                    32'h8b1f03e0,
                    32'h8b1f03e1,
                    32'h8b1f03e2,
                    32'h8b1f03e3,
                    32'h8b040000,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'hd37f3c00,
                    32'h8b040021,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'hd37f3c21,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'h8b080021,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'hf8400022,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'hf8000008,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'hb4fffeff,
                    32'h8b1f03ff,
                    32'h8b1f03ff,
                    32'h8b1f03ff
                };
        
	end
	always_comb begin
		q = ROM[addr];
	end

endmodule


